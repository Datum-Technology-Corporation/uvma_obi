// Copyright 2021 Datum Technology Corporation
// Copyright 2021 Silicon Labs
// Copyright 2021 OpenHW Group
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
// Licensed under the Solderpad Hardware License v 2.1 (the "License"); you may not use this file except in compliance
// with the License, or, at your option, the Apache License version 2.0.  You may obtain a copy of the License at
//                                        https://solderpad.org/licenses/SHL-2.1/
// Unless required by applicable law or agreed to in writing, any work distributed under the License is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.  See the License for the
// specific language governing permissions and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVMT_OBI_ST_DUT_CHKR_SV__
`define __UVMT_OBI_ST_DUT_CHKR_SV__


/**
 * Module encapsulating assertions for Open Bus Interface Agent Self-Testing DUT wrapper (uvmt_obi_st_dut_wrap).
 */
module uvmt_obi_st_dut_chkr(
   uvma_obi_if  mstr_if,
   uvma_obi_if  slv_if
);
   
   // TODO Add assertions to uvmt_obi_st_dut_chkr
   
endmodule : uvmt_obi_st_dut_chkr


`endif // __UVMT_OBI_ST_DUT_CHKR_SV__
