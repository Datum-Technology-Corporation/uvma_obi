// Copyright 2021 Datum Technology Corporation
// Copyright 2021 Silicon Labs
// Copyright 2021 OpenHW Group
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
// Licensed under the Solderpad Hardware License v 2.1 (the "License"); you may not use this file except in compliance
// with the License, or, at your option, the Apache License version 2.0.  You may obtain a copy of the License at
//                                        https://solderpad.org/licenses/SHL-2.1/
// Unless required by applicable law or agreed to in writing, any work distributed under the License is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.  See the License for the
// specific language governing permissions and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_OBI_ST_CHKR_SV__
`define __UVME_OBI_ST_CHKR_SV__


/**
 * TODO Describe uvme_obi_st_chkr
 */
module uvme_obi_st_chkr (
      uvma_obi_if  mstr_if,
      uvma_obi_if  slv_if
);
   
   // TODO Add assertions to uvme_obi_st_chkr
   
endmodule : uvme_obi_st_chkr


`endif // __UVME_OBI_ST_CHKR_SV__
